module reg_group(input clk,we,
input [1:0]raa,
input [1:0]rwba,
input [7:0]i,
output reg[7:0]s,output reg[7:0]d);
reg[7:0] A=8'b0000_0001,B=8'b0000_0010,C=8'b10000000;
parameter a=2'b00,b=2'b01,c=2'b10;

always @(raa or rwba or A or B or C)begin
    
    case (raa)
    a:begin s=A;end
    b:begin s=B;end
    c:begin s=C;end
    default:begin s=1'bz;end
    endcase
    
    case(rwba)
    a:begin d=A;end
    b:begin d=B;end
    c:begin d=C;end
    default:begin d=1'bz;end
    endcase
end

always @(negedge clk)begin

   if(we==1'b0)begin
		if(rwba==a)A<=i;
		else if(rwba==b)B<=i;
		else if(rwba==c)C<=i;
		else A<=A;
    end
    else A<=A;
    
end
endmodule